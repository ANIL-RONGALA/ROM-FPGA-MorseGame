// ECE6370
// Author: ANIL RONGALA, 3848
// My7seg
// This module takes a number as input and produces a 7 bit binary number as an output to control the seven segment display. 


module My7seg(num_input, num_output);
   
   input [3:0] num_input; 
   output [6:0] num_output; 
   reg [6:0] num_output; 

   always @ (num_input)
      begin
         case(num_input)
            4'b0000: begin num_output = 7'b1000000 ; end
            4'b0001: begin num_output = 7'b1111001 ; end
            4'b0010: begin num_output = 7'b0100100 ; end
            4'b0011: begin num_output = 7'b0110000 ; end
            4'b0100: begin num_output = 7'b0011001 ; end
            4'b0101: begin num_output = 7'b0010010 ; end
            4'b0110: begin num_output = 7'b0000010 ; end
            4'b0111: begin num_output = 7'b1111000 ; end
            4'b1000: begin num_output = 7'b0000000 ; end
            4'b1001: begin num_output = 7'b0011000 ; end
            4'b1010: begin num_output = 7'b0001000 ; end 
            4'b1011: begin num_output = 7'b0000011 ; end
            4'b1100: begin num_output = 7'b1000110 ; end
            4'b1101: begin num_output = 7'b0100001 ; end
            4'b1110: begin num_output = 7'b0000110 ; end
            4'b1111: begin num_output = 7'b0001110 ; end
            default: begin num_output = 7'b1111111 ; end
         endcase
      end
endmodule





